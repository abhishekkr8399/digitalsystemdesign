module xor_gate(a, b, y);
 input a;
 input b;
 output y;
 xor G1(y,a,b);
endmodule