module or_gate(a, b, y);
 input a;
 input b;
 output y;
 or G1(y,a,b);
endmodule
