module nor_gate(a, b, y);
 input a;
 input b;
 output y;
 nor G1(y,a,b);
endmodule