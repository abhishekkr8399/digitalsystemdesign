module not_gate(a, y);
 input a;
 output y;
 not G1(y,a);
endmodule
