module and_gate(a, b, y);
 input a;
 input b;
 output y;
 and G1(y,a,b);
endmodule
